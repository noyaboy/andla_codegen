`ifdef ANDLA_CONFIG_VH
`else
`define ANDLA_CONFIG_VH

`define ANDLA_FME_DTYPE "s16"
`define ANDLA_GEMM_I 8
`define ANDLA_IBMC_DATA_BITWIDTH 64
`define ANDLA_GEMM_P 8
`define ANDLA_EDP_E 8
`define ANDLA_BLK_BIU_DATA_WIDTH 64
`define ANDLA_BANK_SIZE 32768
`define ANDLA_IBMC_ADDR_BITWIDTH 19
`define ANDLA_SLV_NUM 16
`define ANDLA_SLV_NUM_BITWIDTH 4
`define ANDLA_SLV0_SUPPORT
`define ANDLA_SLV1_SUPPORT
`define ANDLA_SLV2_SUPPORT
`define ANDLA_SLV3_SUPPORT
`define ANDLA_SLV4_SUPPORT
`define ANDLA_SLV5_SUPPORT
`define ANDLA_SLV6_SUPPORT
`define ANDLA_SLV7_SUPPORT
`define ANDLA_SLV8_SUPPORT
`define ANDLA_SLV9_SUPPORT
`define ANDLA_SLV10_SUPPORT
`define ANDLA_SLV11_SUPPORT
`define ANDLA_SLV12_SUPPORT
`define ANDLA_SLV13_SUPPORT
`define ANDLA_SLV14_SUPPORT
`define ANDLA_SLV15_SUPPORT
`define ANDLA_SHRAM_SIZE_KB 524288
`define ANDLA_512K_SHRAM
`define ANDLA_LDMA_BUFFER_SIZE 256
`define ANDLA_SDMA_BUFFER_SIZE 256
`define ANDLA_LDMA_CMD_FIFO_DEPTH 16
`define ANDLA_SDMA_CMD_FIFO_DEPTH 16
`define ANDLA_FETCH_FIFO_DEPTH 1024
`define ANDLA_FETCH_FIFO_SIZE 4096
`define ANDLA_BIU_BUS axi
`define ANDLA_BUS_AXI
`define ANDLA_BIU_DATA_WIDTH 64
`define ANDLA_BIU_ADDR_WIDTH 32
`define ANDLA_DDMA_SRAM_BUF_EN 1
`define ANDLA_SDMA_SRAM_BUF
`define ANDLA_LDMA_SRAM_BUF
`define ANDLA_CDMA_SRAM_BUF_EN 1
`define ANDLA_CDMA_SRAM_BUF
`define ANDLA_CSR_ID 10711056
`define ANDLA_CSR_REVISION 37888757
`define ANDLA_LDMA_CKSUM_ENABLE 0
`define ANDLA_SDMA_CKSUM_ENABLE 0
`define ANDLA_DDMA_AHB_BRG 0
`define ANDLA_CDMA_AHB_BRG 1
`define ANDLA_ISSUE_AHB_BRG 1
`define ANDLA_LDMA_AHB_BURST_TYPE_EN 0
`define ANDLA_SDMA_AHB_BURST_TYPE_EN 0
`define ANDLA_CDMA_MAX_BURST_LEN 16
`define ANDLA_CDMA_OUTSTD_DEPTH 32

`endif // ANDLA_CONFIG_VH
