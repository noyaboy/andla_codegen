`ifndef ANDLA_VH
`define ANDLA_VH

`include "andla_config.vh"

`ifdef AE350_CONFIG_VH
    `include "config.inc"
    `ifdef ANDLA_BUS_AXI
        `define ANDLA_AXI_SLVID_WIDTH      (`AE350_AXI_ID_WIDTH + 4)
        `define ANDLA_AXI_MSTID_WIDTH      (`AE350_AXI_ID_WIDTH + 0)
        `define ANDLA_AXI_DATA_WIDTH        `NDS_BIU_DATA_WIDTH
        `define ANDLA_DMA_FIFO_DEPTH                         8
        `define ANDLA_AHB_DATA_WIDTH     `NDS_BIU_DATA_WIDTH
        `define ANDLA_AHB_ADDR_WIDTH     `NDS_BIU_ADDR_WIDTH
        `ifdef PLATFORM_FORCE_4GB_SPACE
            `define ANDLA_AXI_ADDR_WIDTH                             32
        `else
            `define ANDLA_AXI_ADDR_WIDTH    `NDS_BIU_ADDR_WIDTH
        `endif // PLATFORM_FORCE_4GB_SPACE
    `else // NDS_IO_AHB
        `define ANDLA_AXI_SLVID_WIDTH      8
        `define ANDLA_AXI_MSTID_WIDTH      8
        `define ANDLA_DMA_FIFO_DEPTH       8
        `ifdef PLATFORM_FORCE_4GB_SPACE 
            `define ANDLA_AXI_ADDR_WIDTH       32
        `else
            `define ANDLA_AXI_ADDR_WIDTH       32
        `endif // PLATFORM_FORCE_4GB_SPACE
        `define ANDLA_AXI_DATA_WIDTH     64
        `define ANDLA_AHB_DATA_WIDTH     `NDS_BIU_DATA_WIDTH
		`ifndef NDS_BIU_ADDR_WIDTH // For Chiuhuahua environment
        	`define ANDLA_AHB_ADDR_WIDTH     32 //`NDS_BIU_ADDR_WIDTH
		`else
        	`define ANDLA_AHB_ADDR_WIDTH     `NDS_BIU_ADDR_WIDTH
        `endif
    `endif
`else
        `define ANDLA_AXI_SLVID_WIDTH                            8
        `define ANDLA_AXI_MSTID_WIDTH                            4
        `define ANDLA_AXI_DATA_WIDTH                            `ANDLA_BLK_BIU_DATA_WIDTH
        `define ANDLA_DMA_FIFO_DEPTH                         8
        `define ANDLA_AXI_ADDR_WIDTH                            `ANDLA_BIU_ADDR_WIDTH
        `define ANDLA_AHB_DATA_WIDTH     `ANDLA_BLK_BIU_DATA_WIDTH
        `define ANDLA_AHB_ADDR_WIDTH     `ANDLA_BIU_ADDR_WIDTH
`endif // AE350_CONFIG

`define ITEM_ID_NUM                     8

`define ANDLA_MAX_PW                    4
`define ANDLA_MAX_PH                    2
`define ANDLA_DLA_OUTSTANDING_DEPTH     4  // defualt 4
`define ANDLA_DLA_SLV_OUTSTANDING_DEPTH     1 
`define ANDLA_DLA_KERNEL_SIZE_BITWIDTH  4  // defualt 15
`define ANDLA_DLA_IMAGE_SIZE_BITWIDTH   10 // defualt 1023
`define ANDLA_DLA_DATA_BITWIDTH         64 // defualt 8
`define ANDLA_DLA_CACC_DATA_BITWIDTH    40 // defualt 40b
`define ANDLA_DLA_BS_DATA_BITWIDTH      32 // defualt 32b
`define ANDLA_DLA_SC_DATA_BITWIDTH      32 // default 32b
`define ANDLA_DLA_TC_DATA_BITWIDTH      32 // defualt 32b

`define ANDLA_IBMC_OUTSTANDING_DEPTH    2
`define ANDLA_MST_NUM                   6
`define ANDLA_MST_NUM_BITWIDTH          3

//LDMA AR/R SETTING
`define ANDLA_LDMA_AR_PENDING_EN  0
`define ANDLA_LDMA_AR_PIPELINE_EN 1
`define ANDLA_LDMA_R_PENDING_EN   1
`define ANDLA_LDMA_R_PIPELINE_EN  1
//LDMA RAM A SETTING
`define ANDLA_LDMA_RAM_ENG_PENDING_EN  1
`define ANDLA_LDMA_RAM_ENG_PIPELINE_EN 0
`define ANDLA_LDMA_RAM_ENG_D_PENDING_EN  1
`define ANDLA_LDMA_RAM_ENG_D_PIPELINE_EN 1
//SDMA AW/W/B SETTING
`define ANDLA_SDMA_AW_PENDING_EN  0
`define ANDLA_SDMA_AW_PIPELINE_EN 1
`define ANDLA_SDMA_W_PENDING_EN   0
`define ANDLA_SDMA_W_PIPELINE_EN  1
`define ANDLA_SDMA_B_PENDING_EN   0
`define ANDLA_SDMA_B_PIPELINE_EN  0

//DMA DATA BUF
`define ANDLA_DMA_SRAM_BUF_EN 1

//`define ANDLA_CDMA_SRAM_BUF_EN `ANDLA_DMA_SRAM_BUF_EN
`define ANDLA_SDMA_SRAM_BUF_EN `ANDLA_DMA_SRAM_BUF_EN
`define ANDLA_LDMA_SRAM_BUF_EN `ANDLA_DMA_SRAM_BUF_EN

`define ITEMID2BASE(x)  ((x << 5) + `ANDLA_REG_BASE

`define ANDLA_SQR_CDMA_FIFO_DEPTH             8
`define ANDLA_SQR_OUTSTANDING_FIFO_DEPTH      2
`define ANDLA_SQR_OUTSTANDING_BUF_DEPTH       2

`define ANDLA_MEM_BASE_ADDRESS                  `ANDLA_AXI_ADDR_WIDTH'hd000_0000
`define ANDLA_REG_BASE_ADDRESS                  `ANDLA_AXI_ADDR_WIDTH'hde00_0000
`define ANDLA_END_ADDRESS                       `ANDLA_AXI_ADDR_WIDTH'hde00_03ff

`define ANDLA_SQR_CREDIT_BITWIDTH             $clog2(`ANDLA_FETCH_FIFO_DEPTH) + 1
`define ANDLA_SQR_INIT_VALUE                  `ANDLA_SQR_CREDIT_BITWIDTH + 2

`define ANDLA_DISP_FIFO_DEPTH                 1024
`define ANDLA_CMD_BITWIDTH                    32
`define ANDLA_RF_WDATA_BITWIDTH               22
`define ANDLA_RF_RDATA_BITWIDTH               32
`define ANDLA_RF_ADDR_BITWIDTH                8
`define ANDLA_RF_ID_BITWIDTH                  3
`define ANDLA_RF_INDEX_BITWIDTH               5

`define ROR_REG_REVISION_PHY_ADDR        `ANDLA_ROR_BASE_ADDRESS + {{(`ANDLA_AXI_ADDR_WIDTH-`ANDLA_RF_INDEX_BITWIDTH-2){1'd0}},(`ANDLA_RF_INDEX_BITWIDTH'd0 << 2)}
`define ROR_REG_ID_PHY_ADDR              `ANDLA_ROR_BASE_ADDRESS + {{(`ANDLA_AXI_ADDR_WIDTH-`ANDLA_RF_INDEX_BITWIDTH-2){1'd0}},(`ANDLA_RF_INDEX_BITWIDTH'd1 << 2)}
`define ROR_REG_STATUS_PHY_ADDR          `ANDLA_ROR_BASE_ADDRESS + {{(`ANDLA_AXI_ADDR_WIDTH-`ANDLA_RF_INDEX_BITWIDTH-2){1'd0}},(`ANDLA_RF_INDEX_BITWIDTH'd2 << 2)}

// autogen_itemid_start
`define CSR_ID        `ANDLA_RF_ID_BITWIDTH'd0
`define SDMA_ID       `ANDLA_RF_ID_BITWIDTH'd1
`define LDMA_ID       `ANDLA_RF_ID_BITWIDTH'd2
`define FME0_ID       `ANDLA_RF_ID_BITWIDTH'd3
`define RESERVED_4_ID `ANDLA_RF_ID_BITWIDTH'd4
`define RESERVED_5_ID `ANDLA_RF_ID_BITWIDTH'd5
`define LDMA2_ID      `ANDLA_RF_ID_BITWIDTH'd6
`define CDMA_ID       `ANDLA_RF_ID_BITWIDTH'd7
// autogen_itemid_stop

`define GEMM_ID                            `ANDLA_RF_ID_BITWIDTH'd5
`define EDP_ID                             `ANDLA_RF_ID_BITWIDTH'd4

`define ANDLA_RF_DDMA_C_SIZE_BITWIDTH           32
`define ANDLA_RF_DDMA_W_SIZE_BITWIDTH           16
`define ANDLA_RF_DDMA_H_SIZE_BITWIDTH           16
`define ANDLA_RF_DDMA_N_SIZE_BITWIDTH           16
`define ANDLA_RF_DDMA_STRIDE_BITWIDTH           32
`define ANDLA_RF_DDMA_PAD_BITWIDTH              4
`define ANDLA_RF_STATUS_BITWIDTH                22
`define ANDLA_RF_CONTROL_BITWIDTH               22
`define ANDLA_RF_CONST_VALUE_BITWIDTH           9

// autogen_provide_common_h_start
`define MODE_BITWIDTH               22
`define CONST_VALUE_BITWIDTH        18
`define RAM_PADDING_VALUE_BITWIDTH  18
`define DILATED_RATE_BITWIDTH       3
`define PAD_SIZE_BITWIDTH           3
`define IM_SIZE_BITWIDTH            14
`define IC_SIZE_BITWIDTH            14
`define KR_SIZE_BITWIDTH            5
// autogen_provide_common_h_stop

`define KC_SIZE_BITWIDTH 14
`define OCBYTE_SIZE_BITWIDTH 14
`define UBMC_ADDR_BITWIDTH `ANDLA_IBMC_ADDR_BITWIDTH

// autogen_bitwidth_start
`define CSR_ID_BITWIDTH                             32
`define CSR_REVISION_BITWIDTH                       32
`define CSR_STATUS_BITWIDTH                         22
`define CSR_CONTROL_BITWIDTH                        22
`define CSR_CREDIT_BITWIDTH                         11
`define CSR_COUNTER_LSB_BITWIDTH                    22
`define CSR_COUNTER_MSB_BITWIDTH                    10
`define CSR_COUNTER_BITWIDTH                        `CSR_COUNTER_LSB_BITWIDTH+`CSR_COUNTER_MSB_BITWIDTH
`define CSR_COUNTER_MASK_BITWIDTH                   22
`define CSR_EXRAM_BASED_ADDR_0_LSB_BITWIDTH         22
`define CSR_EXRAM_BASED_ADDR_0_MSB_BITWIDTH         10
`define CSR_EXRAM_BASED_ADDR_0_BITWIDTH             `CSR_EXRAM_BASED_ADDR_0_LSB_BITWIDTH+`CSR_EXRAM_BASED_ADDR_0_MSB_BITWIDTH
`define CSR_EXRAM_BASED_ADDR_1_LSB_BITWIDTH         22
`define CSR_EXRAM_BASED_ADDR_1_MSB_BITWIDTH         10
`define CSR_EXRAM_BASED_ADDR_1_BITWIDTH             `CSR_EXRAM_BASED_ADDR_1_LSB_BITWIDTH+`CSR_EXRAM_BASED_ADDR_1_MSB_BITWIDTH
`define CSR_EXRAM_BASED_ADDR_2_LSB_BITWIDTH         22
`define CSR_EXRAM_BASED_ADDR_2_MSB_BITWIDTH         10
`define CSR_EXRAM_BASED_ADDR_2_BITWIDTH             `CSR_EXRAM_BASED_ADDR_2_LSB_BITWIDTH+`CSR_EXRAM_BASED_ADDR_2_MSB_BITWIDTH
`define CSR_EXRAM_BASED_ADDR_3_LSB_BITWIDTH         22
`define CSR_EXRAM_BASED_ADDR_3_MSB_BITWIDTH         10
`define CSR_EXRAM_BASED_ADDR_3_BITWIDTH             `CSR_EXRAM_BASED_ADDR_3_LSB_BITWIDTH+`CSR_EXRAM_BASED_ADDR_3_MSB_BITWIDTH
`define CSR_EXRAM_BASED_ADDR_4_LSB_BITWIDTH         22
`define CSR_EXRAM_BASED_ADDR_4_MSB_BITWIDTH         10
`define CSR_EXRAM_BASED_ADDR_4_BITWIDTH             `CSR_EXRAM_BASED_ADDR_4_LSB_BITWIDTH+`CSR_EXRAM_BASED_ADDR_4_MSB_BITWIDTH
`define CSR_EXRAM_BASED_ADDR_5_LSB_BITWIDTH         22
`define CSR_EXRAM_BASED_ADDR_5_MSB_BITWIDTH         10
`define CSR_EXRAM_BASED_ADDR_5_BITWIDTH             `CSR_EXRAM_BASED_ADDR_5_LSB_BITWIDTH+`CSR_EXRAM_BASED_ADDR_5_MSB_BITWIDTH
`define CSR_EXRAM_BASED_ADDR_6_LSB_BITWIDTH         22
`define CSR_EXRAM_BASED_ADDR_6_MSB_BITWIDTH         10
`define CSR_EXRAM_BASED_ADDR_6_BITWIDTH             `CSR_EXRAM_BASED_ADDR_6_LSB_BITWIDTH+`CSR_EXRAM_BASED_ADDR_6_MSB_BITWIDTH
`define CSR_EXRAM_BASED_ADDR_7_LSB_BITWIDTH         22
`define CSR_EXRAM_BASED_ADDR_7_MSB_BITWIDTH         10
`define CSR_EXRAM_BASED_ADDR_7_BITWIDTH             `CSR_EXRAM_BASED_ADDR_7_LSB_BITWIDTH+`CSR_EXRAM_BASED_ADDR_7_MSB_BITWIDTH
`define CSR_NOP_BITWIDTH                            22
`define SDMA_SFENCE_BITWIDTH                        22
`define SDMA_DIRECTION_BITWIDTH                     1
`define SDMA_EXRAM_ADDR_LSB_BITWIDTH                22
`define SDMA_EXRAM_ADDR_MSB_BITWIDTH                10
`define SDMA_EXRAM_ADDR_BITWIDTH                    `SDMA_EXRAM_ADDR_LSB_BITWIDTH+`SDMA_EXRAM_ADDR_MSB_BITWIDTH
`define SDMA_SHRAM_ADDR_BITWIDTH                    `ANDLA_IBMC_ADDR_BITWIDTH
`define SDMA_EXRAM_C_BITWIDTH                       `ANDLA_IBMC_ADDR_BITWIDTH+1
`define SDMA_EXRAM_W_BITWIDTH                       16
`define SDMA_EXRAM_H_BITWIDTH                       16
`define SDMA_EXRAM_N_BITWIDTH                       16
`define SDMA_EXRAM_STRIDE_W_SIZE_BITWIDTH           22
`define SDMA_EXRAM_STRIDE_H_SIZE_BITWIDTH           22
`define SDMA_EXRAM_STRIDE_N_SIZE_BITWIDTH           22
`define SDMA_SHRAM_C_BITWIDTH                       `ANDLA_IBMC_ADDR_BITWIDTH+1
`define SDMA_SHRAM_W_BITWIDTH                       16
`define SDMA_SHRAM_H_BITWIDTH                       16
`define SDMA_SHRAM_N_BITWIDTH                       16
`define SDMA_SHRAM_PAD_RIGHT_BITWIDTH               4
`define SDMA_SHRAM_PAD_LEFT_BITWIDTH                4
`define SDMA_SHRAM_PAD_UP_BITWIDTH                  4
`define SDMA_SHRAM_PAD_DOWN_BITWIDTH                4
`define SDMA_CONST_VALUE_BITWIDTH                   `CONST_VALUE_BITWIDTH
`define SDMA_CH_NUM_BITWIDTH                        `ANDLA_IBMC_ADDR_BITWIDTH+1
`define SDMA_SDMA_DEPADDING_BY_PASS_BITWIDTH        1
`define SDMA_PRESERVED0_BITWIDTH                    1
`define SDMA_PRESERVED1_BITWIDTH                    1
`define SDMA_PRESERVED2_BITWIDTH                    1
`define SDMA_SDMA_CHSUM_SEL_BITWIDTH                22
`define SDMA_SDMA_CHSUM_DATA_BITWIDTH               32
`define SDMA_SHRAM_STRIDE_W_SIZE_BITWIDTH           `ANDLA_IBMC_ADDR_BITWIDTH
`define SDMA_SHRAM_STRIDE_H_SIZE_BITWIDTH           `ANDLA_IBMC_ADDR_BITWIDTH
`define SDMA_SHRAM_STRIDE_N_SIZE_BITWIDTH           `ANDLA_IBMC_ADDR_BITWIDTH
`define LDMA_SFENCE_BITWIDTH                        22
`define LDMA_DIRECTION_BITWIDTH                     1
`define LDMA_EXRAM_ADDR_LSB_BITWIDTH                22
`define LDMA_EXRAM_ADDR_MSB_BITWIDTH                10
`define LDMA_EXRAM_ADDR_BITWIDTH                    `LDMA_EXRAM_ADDR_LSB_BITWIDTH+`LDMA_EXRAM_ADDR_MSB_BITWIDTH
`define LDMA_SHRAM_ADDR_BITWIDTH                    `ANDLA_IBMC_ADDR_BITWIDTH
`define LDMA_EXRAM_C_BITWIDTH                       `ANDLA_IBMC_ADDR_BITWIDTH+1
`define LDMA_EXRAM_W_BITWIDTH                       16
`define LDMA_EXRAM_H_BITWIDTH                       16
`define LDMA_EXRAM_N_BITWIDTH                       16
`define LDMA_EXRAM_STRIDE_W_SIZE_BITWIDTH           22
`define LDMA_EXRAM_STRIDE_H_SIZE_BITWIDTH           22
`define LDMA_EXRAM_STRIDE_N_SIZE_BITWIDTH           22
`define LDMA_SHRAM_C_BITWIDTH                       `ANDLA_IBMC_ADDR_BITWIDTH+1
`define LDMA_SHRAM_W_BITWIDTH                       16
`define LDMA_SHRAM_H_BITWIDTH                       16
`define LDMA_SHRAM_N_BITWIDTH                       16
`define LDMA_SHRAM_PAD_RIGHT_BITWIDTH               4
`define LDMA_SHRAM_PAD_LEFT_BITWIDTH                4
`define LDMA_SHRAM_PAD_UP_BITWIDTH                  4
`define LDMA_SHRAM_PAD_DOWN_BITWIDTH                4
`define LDMA_CONST_VALUE_BITWIDTH                   `CONST_VALUE_BITWIDTH
`define LDMA_CH_NUM_BITWIDTH                        `ANDLA_IBMC_ADDR_BITWIDTH+1
`define LDMA_LDMA_DECOMP_PADDING_BY_PASS_BITWIDTH   1
`define LDMA_RAM_PADDING_VALUE_BITWIDTH             `RAM_PADDING_VALUE_BITWIDTH
`define LDMA_PAD_C_FRONT_BITWIDTH                   14
`define LDMA_PAD_C_BACK_BITWIDTH                    14
`define LDMA_LDMA_CHSUM_SEL_BITWIDTH                22
`define LDMA_LDMA_CHSUM_DATA_BITWIDTH               32
`define LDMA_SHRAM_STRIDE_W_SIZE_BITWIDTH           `ANDLA_IBMC_ADDR_BITWIDTH
`define LDMA_SHRAM_STRIDE_H_SIZE_BITWIDTH           `ANDLA_IBMC_ADDR_BITWIDTH
`define LDMA_SHRAM_STRIDE_N_SIZE_BITWIDTH           `ANDLA_IBMC_ADDR_BITWIDTH
`define FME0_SFENCE_BITWIDTH                        22
`define FME0_MODE_BITWIDTH                          `MODE_BITWIDTH
`define FME0_IM_PAD_BITWIDTH                        `PAD_SIZE_BITWIDTH*4
`define FME0_IM_IW_BITWIDTH                         `IM_SIZE_BITWIDTH
`define FME0_IM_IH_BITWIDTH                         `IM_SIZE_BITWIDTH
`define FME0_IM_IC_BITWIDTH                         `IC_SIZE_BITWIDTH
`define FME0_IM_STRIDE_BITWIDTH                     `KR_SIZE_BITWIDTH*2+4
`define FME0_IM_KERNEL_BITWIDTH                     `KR_SIZE_BITWIDTH*4
`define FME0_OM_OW_BITWIDTH                         `IM_SIZE_BITWIDTH
`define FME0_OM_OH_BITWIDTH                         `IM_SIZE_BITWIDTH
`define FME0_OM_OC_BITWIDTH                         `IC_SIZE_BITWIDTH
`define FME0_IM_ADDR_INIT_BITWIDTH                  `ANDLA_IBMC_ADDR_BITWIDTH
`define FME0_KR_ADDR_INIT_BITWIDTH                  `ANDLA_IBMC_ADDR_BITWIDTH
`define FME0_BS_ADDR_INIT_BITWIDTH                  `ANDLA_IBMC_ADDR_BITWIDTH
`define FME0_PL_ADDR_INIT_BITWIDTH                  `ANDLA_IBMC_ADDR_BITWIDTH
`define FME0_EM_ADDR_INIT_BITWIDTH                  `ANDLA_IBMC_ADDR_BITWIDTH
`define FME0_OM_ADDR_INIT_BITWIDTH                  `ANDLA_IBMC_ADDR_BITWIDTH
`define FME0_EM_ALIGNMENT_ICIW_BITWIDTH             `ANDLA_IBMC_ADDR_BITWIDTH
`define FME0_OM_ALIGNMENT_OCOW_BITWIDTH             `ANDLA_IBMC_ADDR_BITWIDTH
`define FME0_ALIGNMENT_KCKWKH_BITWIDTH              `ANDLA_IBMC_ADDR_BITWIDTH
`define FME0_ALIGNMENT_KCKW_BITWIDTH                `ANDLA_IBMC_ADDR_BITWIDTH
`define FME0_SC_ADDR_INIT_BITWIDTH                  `ANDLA_IBMC_ADDR_BITWIDTH
`define FME0_SH_ADDR_INIT_BITWIDTH                  `ANDLA_IBMC_ADDR_BITWIDTH
`define LDMA2_MODE_CTRL_BITWIDTH                    1
`define LDMA2_ROLL_IC_IW_W_PAD_SIZE_BITWIDTH        `ANDLA_IBMC_ADDR_BITWIDTH+1
`define LDMA2_ROLL_IC_KW_SIZE_BITWIDTH              $clog2(`ANDLA_GEMM_I)+1
`define LDMA2_ROLL_KR_STRIDE_W_SIZE_BITWIDTH        $clog2(`ANDLA_GEMM_I)+1
`define LDMA2_ROLL_PAD_W_LEFT_W_IC_SIZE_BITWIDTH    $clog2(`ANDLA_GEMM_I)+3
`define LDMA2_ROLL_PAD_W_RIGHT_W_IC_SIZE_BITWIDTH   $clog2(`ANDLA_GEMM_I)+3
`define LDMA2_ROLL_PAD_H_SIZE_BITWIDTH              6
`define CDMA_SFENCE_BITWIDTH                        22
`define CDMA_DIRECTION_BITWIDTH                     1
`define CDMA_EXRAM_ADDR_LSB_BITWIDTH                22
`define CDMA_EXRAM_ADDR_MSB_BITWIDTH                10
`define CDMA_EXRAM_ADDR_BITWIDTH                    `CDMA_EXRAM_ADDR_LSB_BITWIDTH+`CDMA_EXRAM_ADDR_MSB_BITWIDTH
`define CDMA_EXRAM_C_BITWIDTH                       22
`define CDMA_EXRAM_W_BITWIDTH                       16
`define CDMA_EXRAM_STRIDE_W_BITWIDTH                22
// autogen_bitwidth_stop

// autogen_idx_start
`define CSR_ID_IDX                            `ANDLA_RF_INDEX_BITWIDTH'd0
`define CSR_REVISION_IDX                      `ANDLA_RF_INDEX_BITWIDTH'd1
`define CSR_STATUS_IDX                        `ANDLA_RF_INDEX_BITWIDTH'd2
`define CSR_CONTROL_IDX                       `ANDLA_RF_INDEX_BITWIDTH'd3
`define CSR_CREDIT_IDX                        `ANDLA_RF_INDEX_BITWIDTH'd4
`define CSR_COUNTER_LSB_IDX                   `ANDLA_RF_INDEX_BITWIDTH'd5
`define CSR_COUNTER_MSB_IDX                   `ANDLA_RF_INDEX_BITWIDTH'd6
`define CSR_COUNTER_MASK_IDX                  `ANDLA_RF_INDEX_BITWIDTH'd7
`define CSR_EXRAM_BASED_ADDR_0_LSB_IDX        `ANDLA_RF_INDEX_BITWIDTH'd8
`define CSR_EXRAM_BASED_ADDR_0_MSB_IDX        `ANDLA_RF_INDEX_BITWIDTH'd9
`define CSR_EXRAM_BASED_ADDR_1_LSB_IDX        `ANDLA_RF_INDEX_BITWIDTH'd10
`define CSR_EXRAM_BASED_ADDR_1_MSB_IDX        `ANDLA_RF_INDEX_BITWIDTH'd11
`define CSR_EXRAM_BASED_ADDR_2_LSB_IDX        `ANDLA_RF_INDEX_BITWIDTH'd12
`define CSR_EXRAM_BASED_ADDR_2_MSB_IDX        `ANDLA_RF_INDEX_BITWIDTH'd13
`define CSR_EXRAM_BASED_ADDR_3_LSB_IDX        `ANDLA_RF_INDEX_BITWIDTH'd14
`define CSR_EXRAM_BASED_ADDR_3_MSB_IDX        `ANDLA_RF_INDEX_BITWIDTH'd15
`define CSR_EXRAM_BASED_ADDR_4_LSB_IDX        `ANDLA_RF_INDEX_BITWIDTH'd16
`define CSR_EXRAM_BASED_ADDR_4_MSB_IDX        `ANDLA_RF_INDEX_BITWIDTH'd17
`define CSR_EXRAM_BASED_ADDR_5_LSB_IDX        `ANDLA_RF_INDEX_BITWIDTH'd18
`define CSR_EXRAM_BASED_ADDR_5_MSB_IDX        `ANDLA_RF_INDEX_BITWIDTH'd19
`define CSR_EXRAM_BASED_ADDR_6_LSB_IDX        `ANDLA_RF_INDEX_BITWIDTH'd20
`define CSR_EXRAM_BASED_ADDR_6_MSB_IDX        `ANDLA_RF_INDEX_BITWIDTH'd21
`define CSR_EXRAM_BASED_ADDR_7_LSB_IDX        `ANDLA_RF_INDEX_BITWIDTH'd22
`define CSR_EXRAM_BASED_ADDR_7_MSB_IDX        `ANDLA_RF_INDEX_BITWIDTH'd23
`define CSR_NOP_IDX                           `ANDLA_RF_INDEX_BITWIDTH'd31
`define SDMA_SFENCE_IDX                       `ANDLA_RF_INDEX_BITWIDTH'd0
`define SDMA_DIRECTION_IDX                    `ANDLA_RF_INDEX_BITWIDTH'd1
`define SDMA_EXRAM_ADDR_LSB_IDX               `ANDLA_RF_INDEX_BITWIDTH'd2
`define SDMA_EXRAM_ADDR_MSB_IDX               `ANDLA_RF_INDEX_BITWIDTH'd3
`define SDMA_SHRAM_ADDR_IDX                   `ANDLA_RF_INDEX_BITWIDTH'd4
`define SDMA_EXRAM_C_IDX                      `ANDLA_RF_INDEX_BITWIDTH'd5
`define SDMA_EXRAM_W_IDX                      `ANDLA_RF_INDEX_BITWIDTH'd6
`define SDMA_EXRAM_H_IDX                      `ANDLA_RF_INDEX_BITWIDTH'd7
`define SDMA_EXRAM_N_IDX                      `ANDLA_RF_INDEX_BITWIDTH'd8
`define SDMA_EXRAM_STRIDE_W_SIZE_IDX          `ANDLA_RF_INDEX_BITWIDTH'd9
`define SDMA_EXRAM_STRIDE_H_SIZE_IDX          `ANDLA_RF_INDEX_BITWIDTH'd10
`define SDMA_EXRAM_STRIDE_N_SIZE_IDX          `ANDLA_RF_INDEX_BITWIDTH'd11
`define SDMA_SHRAM_C_IDX                      `ANDLA_RF_INDEX_BITWIDTH'd12
`define SDMA_SHRAM_W_IDX                      `ANDLA_RF_INDEX_BITWIDTH'd13
`define SDMA_SHRAM_H_IDX                      `ANDLA_RF_INDEX_BITWIDTH'd14
`define SDMA_SHRAM_N_IDX                      `ANDLA_RF_INDEX_BITWIDTH'd15
`define SDMA_SHRAM_PAD_RIGHT_IDX              `ANDLA_RF_INDEX_BITWIDTH'd16
`define SDMA_SHRAM_PAD_LEFT_IDX               `ANDLA_RF_INDEX_BITWIDTH'd17
`define SDMA_SHRAM_PAD_UP_IDX                 `ANDLA_RF_INDEX_BITWIDTH'd18
`define SDMA_SHRAM_PAD_DOWN_IDX               `ANDLA_RF_INDEX_BITWIDTH'd19
`define SDMA_CONST_VALUE_IDX                  `ANDLA_RF_INDEX_BITWIDTH'd20
`define SDMA_CH_NUM_IDX                       `ANDLA_RF_INDEX_BITWIDTH'd21
`define SDMA_SDMA_DEPADDING_BY_PASS_IDX       `ANDLA_RF_INDEX_BITWIDTH'd22
`define SDMA_PRESERVED0_IDX                   `ANDLA_RF_INDEX_BITWIDTH'd23
`define SDMA_PRESERVED1_IDX                   `ANDLA_RF_INDEX_BITWIDTH'd24
`define SDMA_PRESERVED2_IDX                   `ANDLA_RF_INDEX_BITWIDTH'd25
`define SDMA_SDMA_CHSUM_SEL_IDX               `ANDLA_RF_INDEX_BITWIDTH'd26
`define SDMA_SDMA_CHSUM_DATA_IDX              `ANDLA_RF_INDEX_BITWIDTH'd27
`define SDMA_SHRAM_STRIDE_W_SIZE_IDX          `ANDLA_RF_INDEX_BITWIDTH'd28
`define SDMA_SHRAM_STRIDE_H_SIZE_IDX          `ANDLA_RF_INDEX_BITWIDTH'd29
`define SDMA_SHRAM_STRIDE_N_SIZE_IDX          `ANDLA_RF_INDEX_BITWIDTH'd30
`define LDMA_SFENCE_IDX                       `ANDLA_RF_INDEX_BITWIDTH'd0
`define LDMA_DIRECTION_IDX                    `ANDLA_RF_INDEX_BITWIDTH'd1
`define LDMA_EXRAM_ADDR_LSB_IDX               `ANDLA_RF_INDEX_BITWIDTH'd2
`define LDMA_EXRAM_ADDR_MSB_IDX               `ANDLA_RF_INDEX_BITWIDTH'd3
`define LDMA_SHRAM_ADDR_IDX                   `ANDLA_RF_INDEX_BITWIDTH'd4
`define LDMA_EXRAM_C_IDX                      `ANDLA_RF_INDEX_BITWIDTH'd5
`define LDMA_EXRAM_W_IDX                      `ANDLA_RF_INDEX_BITWIDTH'd6
`define LDMA_EXRAM_H_IDX                      `ANDLA_RF_INDEX_BITWIDTH'd7
`define LDMA_EXRAM_N_IDX                      `ANDLA_RF_INDEX_BITWIDTH'd8
`define LDMA_EXRAM_STRIDE_W_SIZE_IDX          `ANDLA_RF_INDEX_BITWIDTH'd9
`define LDMA_EXRAM_STRIDE_H_SIZE_IDX          `ANDLA_RF_INDEX_BITWIDTH'd10
`define LDMA_EXRAM_STRIDE_N_SIZE_IDX          `ANDLA_RF_INDEX_BITWIDTH'd11
`define LDMA_SHRAM_C_IDX                      `ANDLA_RF_INDEX_BITWIDTH'd12
`define LDMA_SHRAM_W_IDX                      `ANDLA_RF_INDEX_BITWIDTH'd13
`define LDMA_SHRAM_H_IDX                      `ANDLA_RF_INDEX_BITWIDTH'd14
`define LDMA_SHRAM_N_IDX                      `ANDLA_RF_INDEX_BITWIDTH'd15
`define LDMA_SHRAM_PAD_RIGHT_IDX              `ANDLA_RF_INDEX_BITWIDTH'd16
`define LDMA_SHRAM_PAD_LEFT_IDX               `ANDLA_RF_INDEX_BITWIDTH'd17
`define LDMA_SHRAM_PAD_UP_IDX                 `ANDLA_RF_INDEX_BITWIDTH'd18
`define LDMA_SHRAM_PAD_DOWN_IDX               `ANDLA_RF_INDEX_BITWIDTH'd19
`define LDMA_CONST_VALUE_IDX                  `ANDLA_RF_INDEX_BITWIDTH'd20
`define LDMA_CH_NUM_IDX                       `ANDLA_RF_INDEX_BITWIDTH'd21
`define LDMA_LDMA_DECOMP_PADDING_BY_PASS_IDX  `ANDLA_RF_INDEX_BITWIDTH'd22
`define LDMA_RAM_PADDING_VALUE_IDX            `ANDLA_RF_INDEX_BITWIDTH'd23
`define LDMA_PAD_C_FRONT_IDX                  `ANDLA_RF_INDEX_BITWIDTH'd24
`define LDMA_PAD_C_BACK_IDX                   `ANDLA_RF_INDEX_BITWIDTH'd25
`define LDMA_LDMA_CHSUM_SEL_IDX               `ANDLA_RF_INDEX_BITWIDTH'd26
`define LDMA_LDMA_CHSUM_DATA_IDX              `ANDLA_RF_INDEX_BITWIDTH'd27
`define LDMA_SHRAM_STRIDE_W_SIZE_IDX          `ANDLA_RF_INDEX_BITWIDTH'd28
`define LDMA_SHRAM_STRIDE_H_SIZE_IDX          `ANDLA_RF_INDEX_BITWIDTH'd29
`define LDMA_SHRAM_STRIDE_N_SIZE_IDX          `ANDLA_RF_INDEX_BITWIDTH'd30
`define FME0_SFENCE_IDX                       `ANDLA_RF_INDEX_BITWIDTH'd0
`define FME0_MODE_IDX                         `ANDLA_RF_INDEX_BITWIDTH'd1
`define FME0_IM_PAD_IDX                       `ANDLA_RF_INDEX_BITWIDTH'd3
`define FME0_IM_IW_IDX                        `ANDLA_RF_INDEX_BITWIDTH'd4
`define FME0_IM_IH_IDX                        `ANDLA_RF_INDEX_BITWIDTH'd5
`define FME0_IM_IC_IDX                        `ANDLA_RF_INDEX_BITWIDTH'd6
`define FME0_IM_STRIDE_IDX                    `ANDLA_RF_INDEX_BITWIDTH'd7
`define FME0_IM_KERNEL_IDX                    `ANDLA_RF_INDEX_BITWIDTH'd8
`define FME0_OM_OW_IDX                        `ANDLA_RF_INDEX_BITWIDTH'd13
`define FME0_OM_OH_IDX                        `ANDLA_RF_INDEX_BITWIDTH'd14
`define FME0_OM_OC_IDX                        `ANDLA_RF_INDEX_BITWIDTH'd15
`define FME0_IM_ADDR_INIT_IDX                 `ANDLA_RF_INDEX_BITWIDTH'd16
`define FME0_KR_ADDR_INIT_IDX                 `ANDLA_RF_INDEX_BITWIDTH'd17
`define FME0_BS_ADDR_INIT_IDX                 `ANDLA_RF_INDEX_BITWIDTH'd18
`define FME0_PL_ADDR_INIT_IDX                 `ANDLA_RF_INDEX_BITWIDTH'd19
`define FME0_EM_ADDR_INIT_IDX                 `ANDLA_RF_INDEX_BITWIDTH'd20
`define FME0_OM_ADDR_INIT_IDX                 `ANDLA_RF_INDEX_BITWIDTH'd21
`define FME0_EM_ALIGNMENT_ICIW_IDX            `ANDLA_RF_INDEX_BITWIDTH'd22
`define FME0_OM_ALIGNMENT_OCOW_IDX            `ANDLA_RF_INDEX_BITWIDTH'd23
`define FME0_ALIGNMENT_KCKWKH_IDX             `ANDLA_RF_INDEX_BITWIDTH'd24
`define FME0_ALIGNMENT_KCKW_IDX               `ANDLA_RF_INDEX_BITWIDTH'd25
`define FME0_SC_ADDR_INIT_IDX                 `ANDLA_RF_INDEX_BITWIDTH'd26
`define FME0_SH_ADDR_INIT_IDX                 `ANDLA_RF_INDEX_BITWIDTH'd27
`define LDMA2_MODE_CTRL_IDX                   `ANDLA_RF_INDEX_BITWIDTH'd0
`define LDMA2_ROLL_IC_IW_W_PAD_SIZE_IDX       `ANDLA_RF_INDEX_BITWIDTH'd1
`define LDMA2_ROLL_IC_KW_SIZE_IDX             `ANDLA_RF_INDEX_BITWIDTH'd2
`define LDMA2_ROLL_KR_STRIDE_W_SIZE_IDX       `ANDLA_RF_INDEX_BITWIDTH'd3
`define LDMA2_ROLL_PAD_W_LEFT_W_IC_SIZE_IDX   `ANDLA_RF_INDEX_BITWIDTH'd4
`define LDMA2_ROLL_PAD_W_RIGHT_W_IC_SIZE_IDX  `ANDLA_RF_INDEX_BITWIDTH'd5
`define LDMA2_ROLL_PAD_H_SIZE_IDX             `ANDLA_RF_INDEX_BITWIDTH'd6
`define CDMA_SFENCE_IDX                       `ANDLA_RF_INDEX_BITWIDTH'd0
`define CDMA_DIRECTION_IDX                    `ANDLA_RF_INDEX_BITWIDTH'd1
`define CDMA_EXRAM_ADDR_LSB_IDX               `ANDLA_RF_INDEX_BITWIDTH'd2
`define CDMA_EXRAM_ADDR_MSB_IDX               `ANDLA_RF_INDEX_BITWIDTH'd3
`define CDMA_EXRAM_C_IDX                      `ANDLA_RF_INDEX_BITWIDTH'd4
`define CDMA_EXRAM_W_IDX                      `ANDLA_RF_INDEX_BITWIDTH'd5
`define CDMA_EXRAM_STRIDE_W_IDX               `ANDLA_RF_INDEX_BITWIDTH'd6
// autogen_idx_stop


`ifdef ANDLA_4M_SHRAM
    `define ANDLA_DLA_CHANNEL_SIZE_BITWIDTH `ANDLA_IBMC_ADDR_BITWIDTH
    `define LDMA_EXRAM_C_BITWIDTH           `UBMC_ADDR_BITWIDTH
    `define LDMA_SHRAM_C_BITWIDTH           `UBMC_ADDR_BITWIDTH
    `define LDMA_CH_NUM_BITWIDTH            `UBMC_ADDR_BITWIDTH
    `define SDMA_EXRAM_C_BITWIDTH           `UBMC_ADDR_BITWIDTH
    `define SDMA_SHRAM_C_BITWIDTH           `UBMC_ADDR_BITWIDTH
    `define SDMA_CH_NUM_BITWIDTH            `UBMC_ADDR_BITWIDTH
`else
    `define ANDLA_DLA_CHANNEL_SIZE_BITWIDTH `ANDLA_IBMC_ADDR_BITWIDTH+1
    `define LDMA_EXRAM_C_BITWIDTH           `UBMC_ADDR_BITWIDTH+1
    `define LDMA_SHRAM_C_BITWIDTH           `UBMC_ADDR_BITWIDTH+1
    `define LDMA_CH_NUM_BITWIDTH            `UBMC_ADDR_BITWIDTH+1
    `define SDMA_EXRAM_C_BITWIDTH           `UBMC_ADDR_BITWIDTH+1
    `define SDMA_SHRAM_C_BITWIDTH           `UBMC_ADDR_BITWIDTH+1
    `define SDMA_CH_NUM_BITWIDTH            `UBMC_ADDR_BITWIDTH+1
`endif

`endif
